
module FA(input a,b,cin,
          output c,s);

assign {c,s} = a+b+cin;

endmodule

