
module butterfly_test();

reg clk,rst;
reg CT;
reg [11:0] A,B,W;
wire[11:0] E,O;
wire[11:0] MUL;
wire[11:0] ADD,SUB;

butterfly uut(clk,rst,
              CT,
              A,B,W,
              E,O,
              MUL,
              ADD,SUB);

always #5 clk = ~clk;

initial begin
    clk = 0;
    rst = 0;
    CT  = 0;
    A   = 0;
    B   = 0;
    W   = 0;

    #200;

    rst = 1;

    #50;
    rst = 0;
    #50;

    A=695;  B=1376; W=1692; CT=0; #10; // E: 2700, O: 3120
    A=518;  B=155;  W=2237; CT=0; #10; // E: 2001, O: 1542
    A=495;  B=331;  W=1996; CT=0; #10; // E: 413, O: 551
    A=2617; B=784;  W=2998; CT=0; #10; // E: 36, O: 1242
    A=80;   B=3195; W=2926; CT=0; #10; // E: 3302, O: 156
    A=2729; B=950;  W=1848; CT=0; #10; // E: 175, O: 2599
    A=763;  B=292;  W=780;  CT=0; #10; // E: 2192, O: 595
    A=258;  B=1629; W=816;  CT=0; #10; // E: 2608, O: 3233

    #100;

    A=3147; B=847;  W=1;    CT=1; #10; // E: 665, O: 2300
    A=2677; B=1496; W=821;  CT=1; #10; // E: 2492, O: 2862
    A=1513; B=2332; W=1476; CT=1; #10; // E: 1359, O: 1667
    A=1936; B=340;  W=2388; CT=1; #10; // E: 1580, O: 2292
    A=1558; B=154;  W=2319; CT=1; #10; // E: 2481, O: 635
    A=3227; B=1516; W=2150; CT=1; #10; // E: 207, O: 2918
    A=2686; B=2702; W=2662; CT=1; #10; // E: 1441, O: 602
    A=1662; B=923;  W=939;  CT=1; #10; // E: 2819, O: 505

end

endmodule
