
module intmul(input [11:0] A,B,
              output[23:0] P);

assign P = A*B;

endmodule
