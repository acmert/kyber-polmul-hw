
/*
The designers:

Ahmet Can Mert <ahmetcanmert@sabanciuniv.edu>
Ferhat Yaman <ferhatyaman@sabanciuniv.edu>

To the extent possible under law, the implementer has waived all copyright
and related or neighboring rights to the source code in this file.
http://creativecommons.org/publicdomain/zero/1.0/
*/


module dt0(
    input [7-1:0] t0_0,
    input [8-1:0] t0_1,
    input [8-1:0] t0_2,
    input [7-1:0] t0_3,
    input [7-1:0] t0_4,
    input [5-1:0] t0_5,
    input [6-1:0] t0_6,
    input [4-1:0] t0_7,
    input [9-1:0] t0_8,
    input [6-1:0] t0_9,
    input [8-1:0] t0_10,
    input [2-1:0] t0_11,
    input [1-1:0] t0_13,
    input [1-1:0] t0_14,
    output [15-1:0] s,
    output [15-1:0] c);

// ------------------------------- Connections

    // --------------------- Level 1

    wire [6-1:0] t1_0;
    wire [6-1:0] t1_1;
    wire [6-1:0] t1_2;
    wire [6-1:0] t1_3;
    wire [6-1:0] t1_4;
    wire [6-1:0] t1_5;
    wire [6-1:0] t1_6;
    wire [5-1:0] t1_7;
    wire [6-1:0] t1_8;
    wire [6-1:0] t1_9;
    wire [6-1:0] t1_10;
    wire [4-1:0] t1_11;
    wire [1-1:0] t1_13;
    wire [1-1:0] t1_14;

    // --------------------- Level 2

    wire [4-1:0] t2_0;
    wire [4-1:0] t2_1;
    wire [4-1:0] t2_2;
    wire [4-1:0] t2_3;
    wire [4-1:0] t2_4;
    wire [4-1:0] t2_5;
    wire [4-1:0] t2_6;
    wire [4-1:0] t2_7;
    wire [4-1:0] t2_8;
    wire [4-1:0] t2_9;
    wire [4-1:0] t2_10;
    wire [4-1:0] t2_11;
    wire [1-1:0] t2_12;
    wire [1-1:0] t2_13;
    wire [1-1:0] t2_14;

    // --------------------- Level 3

    wire [3-1:0] t3_0;
    wire [3-1:0] t3_1;
    wire [3-1:0] t3_2;
    wire [3-1:0] t3_3;
    wire [3-1:0] t3_4;
    wire [3-1:0] t3_5;
    wire [3-1:0] t3_6;
    wire [3-1:0] t3_7;
    wire [3-1:0] t3_8;
    wire [3-1:0] t3_9;
    wire [3-1:0] t3_10;
    wire [3-1:0] t3_11;
    wire [2-1:0] t3_12;
    wire [1-1:0] t3_13;
    wire [1-1:0] t3_14;

    // --------------------- Level 4

    wire [2-1:0] t4_0;
    wire [2-1:0] t4_1;
    wire [2-1:0] t4_2;
    wire [2-1:0] t4_3;
    wire [2-1:0] t4_4;
    wire [2-1:0] t4_5;
    wire [2-1:0] t4_6;
    wire [2-1:0] t4_7;
    wire [2-1:0] t4_8;
    wire [2-1:0] t4_9;
    wire [2-1:0] t4_10;
    wire [2-1:0] t4_11;
    wire [2-1:0] t4_12;
    wire [2-1:0] t4_13;
    wire [1-1:0] t4_14;

// ------------------------------- Operations

    // --------------------- Level 1

    HA u000(t0_0[0],t0_0[1],t1_1[0],t1_0[0]);
    assign t1_0[1] = t0_0[2];
    assign t1_0[2] = t0_0[3];
    assign t1_0[3] = t0_0[4];
    assign t1_0[4] = t0_0[5];
    assign t1_0[5] = t0_0[6];
    FA u010(t0_1[0],t0_1[1],t0_1[2],t1_2[0],t1_1[1]);
    HA u011(t0_1[3],t0_1[4],t1_2[1],t1_1[2]);
    assign t1_1[3] = t0_1[5];
    assign t1_1[4] = t0_1[6];
    assign t1_1[5] = t0_1[7];
    FA u020(t0_2[0],t0_2[1],t0_2[2],t1_3[0],t1_2[2]);
    FA u021(t0_2[3],t0_2[4],t0_2[5],t1_3[1],t1_2[3]);
    assign t1_2[4] = t0_2[6];
    assign t1_2[5] = t0_2[7];
    FA u030(t0_3[0],t0_3[1],t0_3[2],t1_4[0],t1_3[2]);
    HA u031(t0_3[3],t0_3[4],t1_4[1],t1_3[3]);
    assign t1_3[4] = t0_3[5];
    assign t1_3[5] = t0_3[6];
    FA u040(t0_4[0],t0_4[1],t0_4[2],t1_5[0],t1_4[2]);
    HA u041(t0_4[3],t0_4[4],t1_5[1],t1_4[3]);
    assign t1_4[4] = t0_4[5];
    assign t1_4[5] = t0_4[6];
    HA u050(t0_5[0],t0_5[1],t1_6[0],t1_5[2]);
    assign t1_5[3] = t0_5[2];
    assign t1_5[4] = t0_5[3];
    assign t1_5[5] = t0_5[4];
    HA u060(t0_6[0],t0_6[1],t1_7[0],t1_6[1]);
    assign t1_6[2] = t0_6[2];
    assign t1_6[3] = t0_6[3];
    assign t1_6[4] = t0_6[4];
    assign t1_6[5] = t0_6[5];
    assign t1_7[1] = t0_7[0];
    assign t1_7[2] = t0_7[1];
    assign t1_7[3] = t0_7[2];
    assign t1_7[4] = t0_7[3];
    FA u080(t0_8[0],t0_8[1],t0_8[2],t1_9[0],t1_8[0]);
    HA u081(t0_8[3],t0_8[4],t1_9[1],t1_8[1]);
    assign t1_8[2] = t0_8[5];
    assign t1_8[3] = t0_8[6];
    assign t1_8[4] = t0_8[7];
    assign t1_8[5] = t0_8[8];
    FA u090(t0_9[0],t0_9[1],t0_9[2],t1_10[0],t1_9[2]);
    assign t1_9[3] = t0_9[3];
    assign t1_9[4] = t0_9[4];
    assign t1_9[5] = t0_9[5];
    FA u0100(t0_10[0],t0_10[1],t0_10[2],t1_11[0],t1_10[1]);
    HA u0101(t0_10[3],t0_10[4],t1_11[1],t1_10[2]);
    assign t1_10[3] = t0_10[5];
    assign t1_10[4] = t0_10[6];
    assign t1_10[5] = t0_10[7];
    assign t1_11[2] = t0_11[0];
    assign t1_11[3] = t0_11[1];
    assign t1_13[0] = t0_13[0];
    assign t1_14[0] = t0_14[0];

    // --------------------- Level 2

    FA u100(t1_0[0],t1_0[1],t1_0[2],t2_1[0],t2_0[0]);
    assign t2_0[1] = t1_0[3];
    assign t2_0[2] = t1_0[4];
    assign t2_0[3] = t1_0[5];
    FA u110(t1_1[0],t1_1[1],t1_1[2],t2_2[0],t2_1[1]);
    HA u111(t1_1[3],t1_1[4],t2_2[1],t2_1[2]);
    assign t2_1[3] = t1_1[5];
    FA u120(t1_2[0],t1_2[1],t1_2[2],t2_3[0],t2_2[2]);
    FA u121(t1_2[3],t1_2[4],t1_2[5],t2_3[1],t2_2[3]);
    FA u130(t1_3[0],t1_3[1],t1_3[2],t2_4[0],t2_3[2]);
    FA u131(t1_3[3],t1_3[4],t1_3[5],t2_4[1],t2_3[3]);
    FA u140(t1_4[0],t1_4[1],t1_4[2],t2_5[0],t2_4[2]);
    FA u141(t1_4[3],t1_4[4],t1_4[5],t2_5[1],t2_4[3]);
    FA u150(t1_5[0],t1_5[1],t1_5[2],t2_6[0],t2_5[2]);
    FA u151(t1_5[3],t1_5[4],t1_5[5],t2_6[1],t2_5[3]);
    FA u160(t1_6[0],t1_6[1],t1_6[2],t2_7[0],t2_6[2]);
    FA u161(t1_6[3],t1_6[4],t1_6[5],t2_7[1],t2_6[3]);
    FA u170(t1_7[0],t1_7[1],t1_7[2],t2_8[0],t2_7[2]);
    HA u171(t1_7[3],t1_7[4],t2_8[1],t2_7[3]);
    FA u180(t1_8[0],t1_8[1],t1_8[2],t2_9[0],t2_8[2]);
    FA u181(t1_8[3],t1_8[4],t1_8[5],t2_9[1],t2_8[3]);
    FA u190(t1_9[0],t1_9[1],t1_9[2],t2_10[0],t2_9[2]);
    FA u191(t1_9[3],t1_9[4],t1_9[5],t2_10[1],t2_9[3]);
    FA u1100(t1_10[0],t1_10[1],t1_10[2],t2_11[0],t2_10[2]);
    FA u1101(t1_10[3],t1_10[4],t1_10[5],t2_11[1],t2_10[3]);
    FA u1110(t1_11[0],t1_11[1],t1_11[2],t2_12[0],t2_11[2]);
    assign t2_11[3] = t1_11[3];
    assign t2_13[0] = t1_13[0];
    assign t2_14[0] = t1_14[0];

    // --------------------- Level 3

    HA u200(t2_0[0],t2_0[1],t3_1[0],t3_0[0]);
    assign t3_0[1] = t2_0[2];
    assign t3_0[2] = t2_0[3];
    FA u210(t2_1[0],t2_1[1],t2_1[2],t3_2[0],t3_1[1]);
    assign t3_1[2] = t2_1[3];
    FA u220(t2_2[0],t2_2[1],t2_2[2],t3_3[0],t3_2[1]);
    assign t3_2[2] = t2_2[3];
    FA u230(t2_3[0],t2_3[1],t2_3[2],t3_4[0],t3_3[1]);
    assign t3_3[2] = t2_3[3];
    FA u240(t2_4[0],t2_4[1],t2_4[2],t3_5[0],t3_4[1]);
    assign t3_4[2] = t2_4[3];
    FA u250(t2_5[0],t2_5[1],t2_5[2],t3_6[0],t3_5[1]);
    assign t3_5[2] = t2_5[3];
    FA u260(t2_6[0],t2_6[1],t2_6[2],t3_7[0],t3_6[1]);
    assign t3_6[2] = t2_6[3];
    FA u270(t2_7[0],t2_7[1],t2_7[2],t3_8[0],t3_7[1]);
    assign t3_7[2] = t2_7[3];
    FA u280(t2_8[0],t2_8[1],t2_8[2],t3_9[0],t3_8[1]);
    assign t3_8[2] = t2_8[3];
    FA u290(t2_9[0],t2_9[1],t2_9[2],t3_10[0],t3_9[1]);
    assign t3_9[2] = t2_9[3];
    FA u2100(t2_10[0],t2_10[1],t2_10[2],t3_11[0],t3_10[1]);
    assign t3_10[2] = t2_10[3];
    FA u2110(t2_11[0],t2_11[1],t2_11[2],t3_12[0],t3_11[1]);
    assign t3_11[2] = t2_11[3];
    assign t3_12[1] = t2_12[0];
    assign t3_13[0] = t2_13[0];
    assign t3_14[0] = t2_14[0];

    // --------------------- Level 4

    HA u300(t3_0[0],t3_0[1],t4_1[0],t4_0[0]);
    assign t4_0[1] = t3_0[2];
    FA u310(t3_1[0],t3_1[1],t3_1[2],t4_2[0],t4_1[1]);
    FA u320(t3_2[0],t3_2[1],t3_2[2],t4_3[0],t4_2[1]);
    FA u330(t3_3[0],t3_3[1],t3_3[2],t4_4[0],t4_3[1]);
    FA u340(t3_4[0],t3_4[1],t3_4[2],t4_5[0],t4_4[1]);
    FA u350(t3_5[0],t3_5[1],t3_5[2],t4_6[0],t4_5[1]);
    FA u360(t3_6[0],t3_6[1],t3_6[2],t4_7[0],t4_6[1]);
    FA u370(t3_7[0],t3_7[1],t3_7[2],t4_8[0],t4_7[1]);
    FA u380(t3_8[0],t3_8[1],t3_8[2],t4_9[0],t4_8[1]);
    FA u390(t3_9[0],t3_9[1],t3_9[2],t4_10[0],t4_9[1]);
    FA u3100(t3_10[0],t3_10[1],t3_10[2],t4_11[0],t4_10[1]);
    FA u3110(t3_11[0],t3_11[1],t3_11[2],t4_12[0],t4_11[1]);
    HA u3120(t3_12[0],t3_12[1],t4_13[0],t4_12[1]);
    assign t4_13[1] = t3_13[0];
    assign t4_14[0] = t3_14[0];

    // --------------------- Rewire

    assign c[0] = t4_0[0];
    assign c[1] = t4_1[0];
    assign c[2] = t4_2[0];
    assign c[3] = t4_3[0];
    assign c[4] = t4_4[0];
    assign c[5] = t4_5[0];
    assign c[6] = t4_6[0];
    assign c[7] = t4_7[0];
    assign c[8] = t4_8[0];
    assign c[9] = t4_9[0];
    assign c[10] = t4_10[0];
    assign c[11] = t4_11[0];
    assign c[12] = t4_12[0];
    assign c[13] = t4_13[0];
    assign c[14] = t4_14[0];
    assign s[0] = t4_0[1];
    assign s[1] = t4_1[1];
    assign s[2] = t4_2[1];
    assign s[3] = t4_3[1];
    assign s[4] = t4_4[1];
    assign s[5] = t4_5[1];
    assign s[6] = t4_6[1];
    assign s[7] = t4_7[1];
    assign s[8] = t4_8[1];
    assign s[9] = t4_9[1];
    assign s[10] = t4_10[1];
    assign s[11] = t4_11[1];
    assign s[12] = t4_12[1];
    assign s[13] = t4_13[1];
    assign s[14] = 1'b0;

endmodule
